library verilog;
use verilog.vl_types.all;
entity Mux2to1_5bits_tb is
end Mux2to1_5bits_tb;
