library verilog;
use verilog.vl_types.all;
entity Mux4to1_8bits_tb is
end Mux4to1_8bits_tb;
