library verilog;
use verilog.vl_types.all;
entity instructionCycleOp_tb is
end instructionCycleOp_tb;
