library verilog;
use verilog.vl_types.all;
entity Register_5bits_tb is
end Register_5bits_tb;
