library verilog;
use verilog.vl_types.all;
entity instructionSetOp_tb is
end instructionSetOp_tb;
